<?xml version="1.0" encoding="UTF-8"?><Batch version="2.0"><Options AppVersion="7.6.1"><PathAddFiles><![CDATA[C:\Users\arian\OneDrive\Desktop\ariana-portfolio\images\]]></PathAddFiles><PathAddFolder><![CDATA[]]></PathAddFolder></Options><TaskList><Task type="ResizeTask" enabled="true" Comment=""><Width units="0"><![CDATA[960]]></Width><Height units="0"><![CDATA[600]]></Height><DPI><![CDATA[-1]]></DPI><Filter>9</Filter><UseProportions>True</UseProportions><ResizeType>0</ResizeType><ProportionsSize>0</ProportionsSize></Task></TaskList></Batch>